
module unsaved (
	clk_clk,
	reset_reset_n,
	mtl_ip_0_mtl_conduit_export,
	mtl_ip_0_conduit_end_export,
	mtl_ip_0_conduit_end_1_export,
	mtl_ip_0_conduit_end_2_export,
	mtl_ip_0_conduit_end_3_export,
	mtl_ip_0_conduit_end_5_export,
	mtl_ip_0_conduit_end_4_export,
	mtl_ip_0_conduit_end_6_export,
	mtl_ip_0_conduit_end_7_export,
	mtl_ip_0_conduit_end_8_export,
	mtl_ip_0_conduit_end_9_export,
	mtl_ip_0_conduit_end_10_export,
	mtl_ip_0_conduit_end_11_export,
	mtl_ip_0_conduit_end_12_export,
	mtl_ip_0_conduit_end_13_export,
	mtl_ip_0_conduit_end_14_export,
	mtl_ip_0_conduit_end_15_export,
	mtl_ip_0_conduit_end_16_export,
	mtl_ip_0_conduit_end_17_export,
	mtl_ip_0_conduit_end_18_export,
	mtl_ip_0_conduit_end_19_export,
	mtl_ip_0_conduit_end_20_export,
	mtl_ip_0_conduit_end_21_export);	

	input		clk_clk;
	input		reset_reset_n;
	inout		mtl_ip_0_mtl_conduit_export;
	output		mtl_ip_0_conduit_end_export;
	output		mtl_ip_0_conduit_end_1_export;
	output		mtl_ip_0_conduit_end_2_export;
	inout		mtl_ip_0_conduit_end_3_export;
	output	[7:0]	mtl_ip_0_conduit_end_5_export;
	input		mtl_ip_0_conduit_end_4_export;
	output	[7:0]	mtl_ip_0_conduit_end_6_export;
	output	[7:0]	mtl_ip_0_conduit_end_7_export;
	output	[12:0]	mtl_ip_0_conduit_end_8_export;
	output	[1:0]	mtl_ip_0_conduit_end_9_export;
	output		mtl_ip_0_conduit_end_10_export;
	output		mtl_ip_0_conduit_end_11_export;
	output		mtl_ip_0_conduit_end_12_export;
	output		mtl_ip_0_conduit_end_13_export;
	inout	[15:0]	mtl_ip_0_conduit_end_14_export;
	output	[1:0]	mtl_ip_0_conduit_end_15_export;
	output		mtl_ip_0_conduit_end_16_export;
	output		mtl_ip_0_conduit_end_17_export;
	input		mtl_ip_0_conduit_end_18_export;
	input		mtl_ip_0_conduit_end_19_export;
	input		mtl_ip_0_conduit_end_20_export;
	output		mtl_ip_0_conduit_end_21_export;
endmodule
